// adaFruit 32x32 LED display driver